module and_1_bit (
    input wire a,
    input wire b,
    output wire s
);

    assign s = a & b;
    
endmodule